-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Tue Nov 29 21:21:36 2016"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY divider IS 
	PORT
	(
		dividend :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		divisor :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		quotient :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END divider;

ARCHITECTURE bdf_type OF divider IS 

COMPONENT div
	PORT(Si : IN STD_LOGIC;
		 M : IN STD_LOGIC;
		 Bi : IN STD_LOGIC;
		 OKi : IN STD_LOGIC;
		 So : OUT STD_LOGIC;
		 Bo : OUT STD_LOGIC;
		 OKo : OUT STD_LOGIC;
		 D : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	quotient_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_0 <= '0';
SYNTHESIZED_WIRE_13 <= '0';
SYNTHESIZED_WIRE_29 <= '0';
SYNTHESIZED_WIRE_31 <= '0';
SYNTHESIZED_WIRE_48 <= '0';
SYNTHESIZED_WIRE_51 <= '0';
SYNTHESIZED_WIRE_54 <= '0';



b2v_inst : div
PORT MAP(Si => divisor(3),
		 M => SYNTHESIZED_WIRE_0,
		 Bi => SYNTHESIZED_WIRE_1,
		 OKi => SYNTHESIZED_WIRE_2,
		 So => SYNTHESIZED_WIRE_4,
		 Bo => SYNTHESIZED_WIRE_3,
		 OKo => SYNTHESIZED_WIRE_33);


SYNTHESIZED_WIRE_2 <= NOT(SYNTHESIZED_WIRE_3);



b2v_inst11 : div
PORT MAP(Si => SYNTHESIZED_WIRE_4,
		 M => SYNTHESIZED_WIRE_5,
		 Bi => SYNTHESIZED_WIRE_6,
		 OKi => SYNTHESIZED_WIRE_7,
		 So => SYNTHESIZED_WIRE_15,
		 Bo => SYNTHESIZED_WIRE_27,
		 OKo => SYNTHESIZED_WIRE_59);


b2v_inst12 : div
PORT MAP(Si => SYNTHESIZED_WIRE_8,
		 M => SYNTHESIZED_WIRE_9,
		 Bi => SYNTHESIZED_WIRE_10,
		 OKi => SYNTHESIZED_WIRE_11,
		 So => SYNTHESIZED_WIRE_23,
		 Bo => SYNTHESIZED_WIRE_58,
		 OKo => SYNTHESIZED_WIRE_14,
		 D => SYNTHESIZED_WIRE_20);


b2v_inst13 : div
PORT MAP(Si => SYNTHESIZED_WIRE_12,
		 M => dividend(2),
		 Bi => SYNTHESIZED_WIRE_13,
		 OKi => SYNTHESIZED_WIRE_14,
		 So => SYNTHESIZED_WIRE_28,
		 Bo => SYNTHESIZED_WIRE_10,
		 OKo => quotient_ALTERA_SYNTHESIZED(2),
		 D => SYNTHESIZED_WIRE_24);



b2v_inst15 : div
PORT MAP(Si => SYNTHESIZED_WIRE_15,
		 M => SYNTHESIZED_WIRE_16,
		 Bi => SYNTHESIZED_WIRE_17,
		 OKi => SYNTHESIZED_WIRE_18,
		 So => SYNTHESIZED_WIRE_35,
		 Bo => SYNTHESIZED_WIRE_34,
		 OKo => SYNTHESIZED_WIRE_22);


b2v_inst16 : div
PORT MAP(Si => SYNTHESIZED_WIRE_19,
		 M => SYNTHESIZED_WIRE_20,
		 Bi => SYNTHESIZED_WIRE_21,
		 OKi => SYNTHESIZED_WIRE_22,
		 So => SYNTHESIZED_WIRE_39,
		 Bo => SYNTHESIZED_WIRE_17,
		 OKo => SYNTHESIZED_WIRE_26,
		 D => SYNTHESIZED_WIRE_36);


b2v_inst17 : div
PORT MAP(Si => SYNTHESIZED_WIRE_23,
		 M => SYNTHESIZED_WIRE_24,
		 Bi => SYNTHESIZED_WIRE_25,
		 OKi => SYNTHESIZED_WIRE_26,
		 So => SYNTHESIZED_WIRE_43,
		 Bo => SYNTHESIZED_WIRE_21,
		 OKo => SYNTHESIZED_WIRE_30,
		 D => SYNTHESIZED_WIRE_40);


SYNTHESIZED_WIRE_7 <= NOT(SYNTHESIZED_WIRE_27);



b2v_inst19 : div
PORT MAP(Si => SYNTHESIZED_WIRE_28,
		 M => dividend(1),
		 Bi => SYNTHESIZED_WIRE_29,
		 OKi => SYNTHESIZED_WIRE_30,
		 So => SYNTHESIZED_WIRE_47,
		 Bo => SYNTHESIZED_WIRE_25,
		 OKo => quotient_ALTERA_SYNTHESIZED(1),
		 D => SYNTHESIZED_WIRE_44);


b2v_inst2 : div
PORT MAP(Si => divisor(2),
		 M => SYNTHESIZED_WIRE_31,
		 Bi => SYNTHESIZED_WIRE_32,
		 OKi => SYNTHESIZED_WIRE_33,
		 So => SYNTHESIZED_WIRE_56,
		 Bo => SYNTHESIZED_WIRE_1,
		 OKo => SYNTHESIZED_WIRE_53,
		 D => SYNTHESIZED_WIRE_5);


SYNTHESIZED_WIRE_18 <= NOT(SYNTHESIZED_WIRE_34);




b2v_inst22 : div
PORT MAP(Si => SYNTHESIZED_WIRE_35,
		 M => SYNTHESIZED_WIRE_36,
		 Bi => SYNTHESIZED_WIRE_37,
		 OKi => SYNTHESIZED_WIRE_38,
		 Bo => SYNTHESIZED_WIRE_50,
		 OKo => SYNTHESIZED_WIRE_42);

b2v_inst23 : div
PORT MAP(Si => SYNTHESIZED_WIRE_39,
		 M => SYNTHESIZED_WIRE_40,
		 Bi => SYNTHESIZED_WIRE_41,
		 OKi => SYNTHESIZED_WIRE_42,
		 Bo => SYNTHESIZED_WIRE_37,
		 OKo => SYNTHESIZED_WIRE_46);

b2v_inst24 : div
PORT MAP(Si => SYNTHESIZED_WIRE_43,
		 M => SYNTHESIZED_WIRE_44,
		 Bi => SYNTHESIZED_WIRE_45,
		 OKi => SYNTHESIZED_WIRE_46,
		 Bo => SYNTHESIZED_WIRE_41,
		 OKo => SYNTHESIZED_WIRE_49);

b2v_inst25 : div
PORT MAP(Si => SYNTHESIZED_WIRE_47,
		 M => dividend(0),
		 Bi => SYNTHESIZED_WIRE_48,
		 OKi => SYNTHESIZED_WIRE_49,
		 Bo => SYNTHESIZED_WIRE_45,
		 OKo => quotient_ALTERA_SYNTHESIZED(0));

SYNTHESIZED_WIRE_38 <= NOT(SYNTHESIZED_WIRE_50);




b2v_inst3 : div
PORT MAP(Si => divisor(1),
		 M => SYNTHESIZED_WIRE_51,
		 Bi => SYNTHESIZED_WIRE_52,
		 OKi => SYNTHESIZED_WIRE_53,
		 So => SYNTHESIZED_WIRE_8,
		 Bo => SYNTHESIZED_WIRE_32,
		 OKo => SYNTHESIZED_WIRE_55,
		 D => SYNTHESIZED_WIRE_57);


b2v_inst4 : div
PORT MAP(Si => divisor(0),
		 M => dividend(3),
		 Bi => SYNTHESIZED_WIRE_54,
		 OKi => SYNTHESIZED_WIRE_55,
		 So => SYNTHESIZED_WIRE_12,
		 Bo => SYNTHESIZED_WIRE_52,
		 OKo => quotient_ALTERA_SYNTHESIZED(3),
		 D => SYNTHESIZED_WIRE_9);


b2v_inst5 : div
PORT MAP(Si => SYNTHESIZED_WIRE_56,
		 M => SYNTHESIZED_WIRE_57,
		 Bi => SYNTHESIZED_WIRE_58,
		 OKi => SYNTHESIZED_WIRE_59,
		 So => SYNTHESIZED_WIRE_19,
		 Bo => SYNTHESIZED_WIRE_6,
		 OKo => SYNTHESIZED_WIRE_11,
		 D => SYNTHESIZED_WIRE_16);





quotient <= quotient_ALTERA_SYNTHESIZED;

END bdf_type;